module and6 (
    input  [5:0] a,
    input  [5:0] b,
    output [5:0] y
);
  assign y = a & b;
endmodule
